`timescale 1 ns/10 ps

`define	TestPort1	30'h0 
`define	TestPort2	30'h1  
`define	TestPort3	30'h2  
`define	TestPort4	30'h3  
`define	TestPort5	30'h4 
`define	TestPort6	30'h5  
`define	TestPort7	30'h6  
`define	TestPort8	30'h7  
`define	TestPort9	30'h8 
`define	TestPort10	30'h9  
`define	TestPort11	30'hA  
`define	TestPort12	30'hB  
`define	TestPort13	30'hC 
`define	TestPort14	30'hD  

`define	answer1	 32'hFFFFFFFE
`define	answer2	 32'h00000002
`define	answer3	 32'h00000007
`define	answer4	 32'h00000001
`define	answer5	 32'hFFFFFFFF
`define	answer6	 32'h00000003
`define	answer7	 32'h00000000
`define	answer8	 32'hFFFFFFFF
`define	answer9	 32'hFFFFFFFF
`define	answer10 32'hFFFFFFFC
`define	answer11 32'h00000001
`define	answer12 32'hFFFFFFFF
`define	answer13 32'h00000000
`define	answer14 32'hFFFFFFFE

`define	CheckNum	6'd13

module	TestBed(
	clk,
	rst,
	addr,
	data,
	wen,
	error_num,
	duration,
	finish
);
	input			clk, rst;
	input	[29:0]	addr;
	input	[31:0]	data;
	input			wen;
	output	[7:0]	error_num;
	output	[15:0]	duration;
	output			finish;
	reg		[7:0]	error_num;
	reg		[15:0]	duration;
	reg				finish;
	
	reg		[1:0]	curstate;
	reg		[1:0]	nxtstate;
	reg		[5:0]	curaddr;
	reg		[5:0]	nxtaddr;
	reg		[15:0]	nxtduration;
	reg		[7:0]	nxt_error_num;
	reg				state,state_next;

	wire     [31:0]  data_modify;
		
	parameter	state_idle 	= 2'b00;
	parameter	state_check= 2'b01;
	parameter	state_report= 2'b10;	
		
	assign data_modify = {data[7:0],data[15:8],data[23:16],data[31:24]}; // convert little-endian format to readable format

	always@( posedge clk or negedge rst )						// State-DFF
	begin
		if( ~rst )
		begin
			curstate <= state_idle;
			curaddr  <= 0;
			duration <= 0;
			error_num <= 8'd255;
			
			state <= 0;
		end
		else
		begin
			curstate <= nxtstate;
			curaddr  <= nxtaddr;
			duration <= nxtduration;
			error_num <= nxt_error_num;
			
			state <= state_next;
		end
	end
			
	always@(negedge clk)	// FSM for test
	begin
		finish = 1'b0;
		case( curstate )
		state_idle: 	begin
							nxtaddr = 0;
							nxtduration = 0;
							nxt_error_num = 255;	
							if( addr==`TestPort1 && data_modify==`answer1 && wen )
							begin
								nxt_error_num = 0;
								nxtstate = state_check;
								nxtaddr = 1;
							end	 	
							else nxtstate = state_idle;
						end
		state_check:	begin
							nxtduration = duration + 1;
							nxtaddr = curaddr;						
							nxt_error_num = error_num;	
							if( addr==`TestPort2 && wen && state==0 )
							begin
								// $display("2: %h %h",data_modify, `answer2);
								nxtaddr = addr + 1; 
								if( data_modify != `answer2 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 2: %h %h",data_modify, `answer2);
								end
							end
							else if( addr==`TestPort3 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer3 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 3: %h %h",data_modify, `answer3);
								end
							end
							else if( addr==`TestPort4 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer4 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 4: %h %h",data_modify, `answer4);
								end
							end
							else if( addr==`TestPort5 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer5 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 5: %h %h",data_modify, `answer5);
								end
							end
							else if( addr==`TestPort6 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer6 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 6: %h %h",data_modify, `answer6);
								end
							end
							else if( addr==`TestPort7 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer7 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 7: %h %h",data_modify, `answer7);
								end
							end
							else if( addr==`TestPort8 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer8 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 8: %h %h",data_modify, `answer8);
								end
							end
							else if( addr==`TestPort9 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer9 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 9: %h %h",data_modify, `answer9);
								end
							end
							else if( addr==`TestPort10 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer10 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 10: %h %h",data_modify, `answer10);
								end
							end
							else if( addr==`TestPort11 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer11 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 11: %h %h",data_modify, `answer11);
								end
							end
							else if( addr==`TestPort12 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer12 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 12: %h %h",data_modify, `answer12);
								end
							end
							else if( addr==`TestPort13 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer13 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 13: %h %h",data_modify, `answer13);
								end
							end
							else if( addr==`TestPort14 && wen && state==0 )
							begin
								nxtaddr = addr + 1;
								if( data_modify != `answer14 ) begin
									nxt_error_num = error_num + 8'd1;
									$display("Error at 14: %h %h",data_modify, `answer14);
								end
							end

							nxtstate = curstate;
							if( addr==`CheckNum )	
								nxtstate = state_report;
						end
		state_report:	begin
							finish = 1'b1;
							nxtaddr = curaddr;
							nxtstate = curstate;		
							nxtduration = duration;
							nxt_error_num = error_num;	
						end						
		endcase	
	end
	
	always@(*)begin//sub-FSM (avoid the Dcache stall condition)
		case(state)
			1'b0:begin
				if(wen)
					state_next=1;
				else
					state_next=state;				
			end
			1'b1:begin
				if(!wen)
					state_next=0;
				else
					state_next=state;	
			end
		endcase
	end

	always@( negedge clk )						
	begin
		if(curstate == state_report) begin
			$display("--------------------------- Simulation FINISH !!---------------------------");
			if (error_num) begin 
				$display("============================================================================");
				$display("\n (T_T) FAIL!! The simulation result is FAIL!!! there were %d errors at all.\n", error_num);
				$display("============================================================================");
			end
			 else begin 
				$display("============================================================================");
				$display("\n \\(^o^)/ CONGRATULATIONS!!  The simulation result is PASS!!!\n");
				$display("============================================================================");
			end
		end
	end
endmodule
